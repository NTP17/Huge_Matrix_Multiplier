module adder17 (
	input [16:0] D, E,
	output [17:0] F
);

	assign F = E + D;

endmodule