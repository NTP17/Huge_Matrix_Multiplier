module multiplier_8816 (
	dataa,
	datab,
	result);

	input	[7:0]  dataa;
	input	[7:0]  datab;
	output	[15:0]  result;

	assign result = dataa * datab;

endmodule