// megafunction wizard: %PARALLEL_ADD%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: parallel_add 

// ============================================================
// File Name: adder18.v
// Megafunction Name(s):
// 			parallel_add
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 18.1.0 Build 625 09/12/2018 SJ Lite Edition
// ************************************************************


//Copyright (C) 2018  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module adder18 (
	data0x,
	data1x,
	data2x,
	data3x,
	data4x,
	data5x,
	data6x,
	data7x,
	data8x,
	result);

	input	[17:0]  data0x;
	input	[17:0]  data1x;
	input	[17:0]  data2x;
	input	[17:0]  data3x;
	input	[17:0]  data4x;
	input	[17:0]  data5x;
	input	[17:0]  data6x;
	input	[17:0]  data7x;
	input	[17:0]  data8x;
	output	[21:0]  result;

	wire [21:0] sub_wire10;
	wire [17:0] sub_wire9 = data8x[17:0];
	wire [17:0] sub_wire8 = data7x[17:0];
	wire [17:0] sub_wire7 = data6x[17:0];
	wire [17:0] sub_wire6 = data5x[17:0];
	wire [17:0] sub_wire5 = data4x[17:0];
	wire [17:0] sub_wire4 = data3x[17:0];
	wire [17:0] sub_wire3 = data2x[17:0];
	wire [17:0] sub_wire2 = data1x[17:0];
	wire [17:0] sub_wire0 = data0x[17:0];
	wire [161:0] sub_wire1 = {sub_wire9, sub_wire8, sub_wire7, sub_wire6, sub_wire5, sub_wire4, sub_wire3, sub_wire2, sub_wire0};
	wire [21:0] result = sub_wire10[21:0];

	parallel_add	parallel_add_component (
				.data (sub_wire1),
				.result (sub_wire10)
				// synopsys translate_off
				,
				.aclr (),
				.clken (),
				.clock ()
				// synopsys translate_on
				);
	defparam
		parallel_add_component.msw_subtract = "NO",
		parallel_add_component.pipeline = 0,
		parallel_add_component.representation = "UNSIGNED",
		parallel_add_component.result_alignment = "LSB",
		parallel_add_component.shift = 0,
		parallel_add_component.size = 9,
		parallel_add_component.width = 18,
		parallel_add_component.widthr = 22;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: MSW_SUBTRACT STRING "NO"
// Retrieval info: CONSTANT: PIPELINE NUMERIC "0"
// Retrieval info: CONSTANT: REPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: RESULT_ALIGNMENT STRING "LSB"
// Retrieval info: CONSTANT: SHIFT NUMERIC "0"
// Retrieval info: CONSTANT: SIZE NUMERIC "9"
// Retrieval info: CONSTANT: WIDTH NUMERIC "18"
// Retrieval info: CONSTANT: WIDTHR NUMERIC "22"
// Retrieval info: USED_PORT: data0x 0 0 18 0 INPUT NODEFVAL "data0x[17..0]"
// Retrieval info: USED_PORT: data1x 0 0 18 0 INPUT NODEFVAL "data1x[17..0]"
// Retrieval info: USED_PORT: data2x 0 0 18 0 INPUT NODEFVAL "data2x[17..0]"
// Retrieval info: USED_PORT: data3x 0 0 18 0 INPUT NODEFVAL "data3x[17..0]"
// Retrieval info: USED_PORT: data4x 0 0 18 0 INPUT NODEFVAL "data4x[17..0]"
// Retrieval info: USED_PORT: data5x 0 0 18 0 INPUT NODEFVAL "data5x[17..0]"
// Retrieval info: USED_PORT: data6x 0 0 18 0 INPUT NODEFVAL "data6x[17..0]"
// Retrieval info: USED_PORT: data7x 0 0 18 0 INPUT NODEFVAL "data7x[17..0]"
// Retrieval info: USED_PORT: data8x 0 0 18 0 INPUT NODEFVAL "data8x[17..0]"
// Retrieval info: USED_PORT: result 0 0 22 0 OUTPUT NODEFVAL "result[21..0]"
// Retrieval info: CONNECT: @data 0 0 18 0 data0x 0 0 18 0
// Retrieval info: CONNECT: @data 0 0 18 18 data1x 0 0 18 0
// Retrieval info: CONNECT: @data 0 0 18 36 data2x 0 0 18 0
// Retrieval info: CONNECT: @data 0 0 18 54 data3x 0 0 18 0
// Retrieval info: CONNECT: @data 0 0 18 72 data4x 0 0 18 0
// Retrieval info: CONNECT: @data 0 0 18 90 data5x 0 0 18 0
// Retrieval info: CONNECT: @data 0 0 18 108 data6x 0 0 18 0
// Retrieval info: CONNECT: @data 0 0 18 126 data7x 0 0 18 0
// Retrieval info: CONNECT: @data 0 0 18 144 data8x 0 0 18 0
// Retrieval info: CONNECT: result 0 0 22 0 @result 0 0 22 0
// Retrieval info: GEN_FILE: TYPE_NORMAL adder18.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL adder18.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL adder18.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL adder18.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL adder18_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL adder18_bb.v FALSE
// Retrieval info: LIB_FILE: altera_mf
